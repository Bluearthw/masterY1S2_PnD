// Digital version of biasing
module biasing (
    output wire vdd,
    output wire vss,
    output wire comp_ref
  );
endmodule

