// Digital version of anatop_driver
module anatop_driver (output wire out);
endmodule
