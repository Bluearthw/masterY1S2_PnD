//Verilog HDL for "PnD", "vga_ctrl_v1" "functional"


module vga_ctrl_v1 ( );

endmodule
